module alu
(
    input logic         clk, 
    input logic[31:0]   a,
    input logic[31:0]   b,
    input logic[1:0]    op,
    output logic[31:0]  res
);

    always @(posedge clk) begin;
        
    end

endmodule