module main();

endmodule