module xor32
(
    input logic[31:0]   i,
    output wire         o
);
    assign o = ^o;

endmodule

module or32
(
    input logic[31:0]   i,
    output wire         o
);
    

endmodule