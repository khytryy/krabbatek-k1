module main;
    initial begin
        $display("Krabba!");
        $finish;
    end
endmodule